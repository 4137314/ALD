# modello BRAM semplice