# array NxN di PE