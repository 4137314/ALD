# Multiply-Accumulate unit