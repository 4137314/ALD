# sequenziatore principale