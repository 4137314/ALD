mat2x2_accel.vhd