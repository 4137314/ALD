# top-level TPU