# Processing Element (1 MAC + activation)